library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b98",x"ad040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b98",x"c9040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"c3040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88a6",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9e",x"a0738306",x"10100508",x"060b0b0b",x"88a90400",x"00000000",x"00000000",x"0b0b0b88",x"f7040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"df040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9ee80c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d43f95",x"ef3f0410",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10105351",x"047381ff",x"06738306",x"09810583",x"05101010",x"2b0772fc",x"060c5151",x"043c0472",x"72807281",x"06ff0509",x"72060571",x"1052720a",x"100a5372",x"ed385151",x"53510488",x"088c0890",x"08757599",x"a22d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"08757598",x"de2d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"088df62d",x"900c8c0c",x"880c04ff",x"3d0d0b0b",x"0b9ef833",x"5170a638",x"9ef40870",x"08525270",x"802e9238",x"84129ef4",x"0c702d9e",x"f4087008",x"525270f0",x"38810b0b",x"0b0b9ef8",x"34833d0d",x"0404803d",x"0d0b0b0b",x"9fa40880",x"2e8e380b",x"0b0b0b80",x"0b802e09",x"81068538",x"823d0d04",x"0b0b0b9f",x"a4510b0b",x"0bf6813f",x"823d0d04",x"04ff3d0d",x"80c48080",x"84527108",x"70822a70",x"81065151",x"5170f338",x"833d0d04",x"ff3d0d80",x"c4808084",x"52710870",x"812a7081",x"06515151",x"70f33873",x"82900a0c",x"833d0d04",x"fe3d0d74",x"7080dc80",x"80880c70",x"81ff06ff",x"83115451",x"53718126",x"8d3880fd",x"518aa02d",x"72a03251",x"83397251",x"8aa02d84",x"3d0d0480",x"3d0d83ff",x"ff0b83d0",x"0a0c80fe",x"518aa02d",x"823d0d04",x"ff3d0d83",x"d00a0870",x"882a5252",x"8ac02d71",x"81ff0651",x"8ac02d80",x"fe518aa0",x"2d833d0d",x"0482f6ff",x"0b80cc80",x"80880c80",x"0b80cc80",x"80840c9f",x"0b83900a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808470",x"08708480",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80847008",x"70fbffff",x"06720c52",x"52833d0d",x"04a0900b",x"a0800c9e",x"fc0ba084",x"0c98c22d",x"ff3d0d73",x"518b710c",x"90115298",x"8080720c",x"80720c70",x"0883ffff",x"06880c83",x"3d0d04fa",x"3d0d787a",x"7dff1e57",x"57585373",x"ff2ea738",x"80568452",x"75730c72",x"0888180c",x"ff125271",x"f3387484",x"16740872",x"0cff1656",x"565273ff",x"2e098106",x"dd38883d",x"0d04f83d",x"0d80d080",x"80845783",x"d00a598b",x"da2d7651",x"8c802d9e",x"fc708808",x"10109880",x"84057170",x"8405530c",x"5656fb80",x"84a1ad75",x"0c9ed80b",x"88170c80",x"70780c77",x"0c760883",x"ffff0656",x"81df800b",x"88082783",x"38ff3983",x"ffff790c",x"a0805488",x"08537852",x"76518c9f",x"2d76518b",x"be2d7808",x"5574762e",x"893880c3",x"518aa02d",x"ff39a084",x"085574fb",x"a0849e80",x"2e893880",x"c2518aa0",x"2dff3980",x"d00a7008",x"70ffbf06",x"720c5656",x"8a852d8b",x"f12dff3d",x"0d9f8808",x"81119f88",x"0c518390",x"0a700870",x"feff0672",x"0c525283",x"3d0d0480",x"3d0d8aef",x"2d728180",x"07518ac0",x"2d8b842d",x"823d0d04",x"fe3d0d80",x"d0808084",x"538bda2d",x"85730c80",x"730c7208",x"7081ff06",x"74535152",x"8bbe2d71",x"880c843d",x"0d04fc3d",x"0d768111",x"33821233",x"7181800a",x"29718480",x"80290583",x"14337082",x"80291284",x"16335271",x"05a08005",x"86168517",x"33575253",x"53555755",x"53ff1353",x"72ff2e91",x"38737081",x"05553352",x"71757081",x"055734e9",x"3989518e",x"932d863d",x"0d04f93d",x"0d795780",x"d0808084",x"568bda2d",x"81173382",x"18337182",x"80290553",x"5371802e",x"94388517",x"72555372",x"70810554",x"33760cff",x"145473f3",x"38831733",x"84183371",x"82802905",x"56528054",x"73752797",x"38735877",x"760c7614",x"76085353",x"71733481",x"14547474",x"26ed3875",x"518bbe2d",x"8aef2d81",x"84518ac0",x"2d74882a",x"518ac02d",x"74518ac0",x"2d805473",x"75278f38",x"76147033",x"52528ac0",x"2d811454",x"ee398b84",x"2d893d0d",x"04f93d0d",x"795680d0",x"80808455",x"8bda2d86",x"750c7451",x"8bbe2d8b",x"da2d81ad",x"70760c81",x"17338218",x"33718280",x"29058319",x"33780c84",x"1933780c",x"85193378",x"0c595353",x"80547377",x"27b33872",x"5873802e",x"87388bda",x"2d77750c",x"73168611",x"33760c87",x"1133760c",x"5274518b",x"be2d8ea8",x"2d880881",x"065271f6",x"38821454",x"767426d1",x"388bda2d",x"84750c74",x"518bbe2d",x"8aef2d81",x"87518ac0",x"2d8b842d",x"893d0d04",x"fc3d0d76",x"81113382",x"12337190",x"2b71882b",x"07831433",x"70720788",x"2b841633",x"71075152",x"53575754",x"5288518e",x"932d81ff",x"518aa02d",x"80c48080",x"84537208",x"70812a70",x"81065151",x"5271f338",x"73848080",x"0780c480",x"80840c86",x"3d0d04fe",x"3d0d8ea8",x"2d880888",x"08810653",x"5371f338",x"8aef2d81",x"83518ac0",x"2d72518a",x"c02d8b84",x"2d843d0d",x"04fe3d0d",x"800b9f88",x"0c8aef2d",x"8181518a",x"c02d9ed8",x"538f5272",x"70810554",x"33518ac0",x"2dff1252",x"71ff2e09",x"8106ec38",x"8b842d84",x"3d0d04fe",x"3d0d800b",x"9f880c8a",x"ef2d8182",x"518ac02d",x"80d08080",x"84528bda",x"2d81f90a",x"0b80d080",x"809c0c71",x"08725253",x"8bbe2d72",x"9f900c72",x"902a518a",x"c02d9f90",x"08882a51",x"8ac02d9f",x"9008518a",x"c02d8ea8",x"2d880851",x"8ac02d8b",x"842d843d",x"0d04803d",x"0d810b9f",x"8c0c800b",x"83900a0c",x"85518e93",x"2d823d0d",x"04803d0d",x"800b9f8c",x"0c8ba52d",x"86518e93",x"2d823d0d",x"04fd3d0d",x"80d08080",x"84548a51",x"8e932d8b",x"da2d9efc",x"7452538c",x"802d7288",x"08101098",x"80840571",x"70840553",x"0c52fb80",x"84a1ad72",x"0c9ed80b",x"88140c73",x"518bbe2d",x"8a852d8b",x"f12dfc3d",x"0d80d080",x"80847052",x"558bbe2d",x"8bda2d8b",x"750c7680",x"d0808094",x"0c80750c",x"a0805477",x"5383d00a",x"5274518c",x"9f2d7451",x"8bbe2d8a",x"852d8bf1",x"2dffab3d",x"0d800b9f",x"8c0c800b",x"9f880c80",x"0b8df60b",x"a0800c57",x"80c48080",x"84558480",x"b3750c80",x"c88080a4",x"53fbffff",x"73087072",x"06750c53",x"5480c880",x"80947008",x"70760672",x"0c5353a8",x"7099da71",x"70840553",x"0c9ab771",x"0c539bd0",x"0b88120c",x"9cdf0b8c",x"120c94b2",x"0b90120c",x"53880b80",x"c0808084",x"0c900a53",x"81730c8b",x"a52dfe88",x"880b80dc",x"8080840c",x"81f20b80",x"d00a0c80",x"d0808084",x"7052528b",x"be2d8bda",x"2d71518b",x"be2d8bda",x"2d84720c",x"71518bbe",x"2d8bda2d",x"86720c71",x"518bbe2d",x"8bda2d81",x"98720c71",x"518bbe2d",x"76777675",x"933d4141",x"5b5b5b83",x"d00a5c78",x"08708106",x"5152719d",x"389f8c08",x"5372f038",x"9f880852",x"87e87227",x"e638727e",x"0c728390",x"0a0c98bb",x"2d82900a",x"08537980",x"2e81b438",x"7280fe2e",x"09810680",x"f4387680",x"2ec13880",x"7d785856",x"5a827727",x"ffb53883",x"ffff7c0c",x"79fe1853",x"53797227",x"983880dc",x"80808872",x"55587413",x"7033790c",x"52811353",x"737326f2",x"38ff1670",x"16547505",x"ff057033",x"74337072",x"882b077f",x"08535155",x"51527173",x"2e098106",x"feed3874",x"3353728a",x"26fee438",x"7210109e",x"ac057552",x"70085152",x"712dfed3",x"397280fd",x"2e098106",x"8638815b",x"fec53976",x"829f269e",x"387a802e",x"87388073",x"a032545b",x"80d73d77",x"05fde005",x"52727234",x"811757fe",x"a239805a",x"fe9d3972",x"80fe2e09",x"8106fe93",x"387957ff",x"7c0c8177",x"5c5afe87",x"39ff3d0d",x"80528051",x"94e92d83",x"3d0d0481",x"fff80d8c",x"da0481ff",x"f80da088",x"04880880",x"c0808088",x"08a08008",x"2d50880c",x"810b900a",x"0c04fb3d",x"0d777955",x"55805675",x"7524ab38",x"8074249d",x"38805373",x"52745180",x"e13f8808",x"5475802e",x"85388808",x"30547388",x"0c873d0d",x"04733076",x"81325754",x"dc397430",x"55815673",x"8025d238",x"ec39fa3d",x"0d787a57",x"55805776",x"7524a438",x"759f2c54",x"81537574",x"32743152",x"74519b3f",x"88085476",x"802e8538",x"88083054",x"73880c88",x"3d0d0474",x"30558157",x"d739fc3d",x"0d767853",x"54815380",x"74732652",x"5572802e",x"98387080",x"2ea93880",x"7224a438",x"71107310",x"75722653",x"545272ea",x"38735178",x"83387451",x"70880c86",x"3d0d0472",x"812a7281",x"2a535372",x"802ee638",x"717426ef",x"38737231",x"75740774",x"812a7481",x"2a555556",x"54e539fc",x"3d0d7670",x"797b5555",x"55558f72",x"278c3872",x"75078306",x"5170802e",x"a738ff12",x"5271ff2e",x"98387270",x"81055433",x"74708105",x"5634ff12",x"5271ff2e",x"098106ea",x"3874880c",x"863d0d04",x"74517270",x"84055408",x"71708405",x"530c7270",x"84055408",x"71708405",x"530c7270",x"84055408",x"71708405",x"530c7270",x"84055408",x"71708405",x"530cf012",x"52718f26",x"c9388372",x"27953872",x"70840554",x"08717084",x"05530cfc",x"12527183",x"26ed3870",x"54ff8339",x"fc3d0d76",x"7971028c",x"059f0533",x"57555355",x"8372278a",x"38748306",x"5170802e",x"a238ff12",x"5271ff2e",x"93387373",x"70810555",x"34ff1252",x"71ff2e09",x"8106ef38",x"74880c86",x"3d0d0474",x"74882b75",x"07707190",x"2b075154",x"518f7227",x"a5387271",x"70840553",x"0c727170",x"8405530c",x"72717084",x"05530c72",x"71708405",x"530cf012",x"52718f26",x"dd388372",x"27903872",x"71708405",x"530cfc12",x"52718326",x"f2387053",x"ff9039fb",x"3d0d7779",x"70720783",x"06535452",x"70933871",x"73730854",x"56547173",x"082e80c4",x"38737554",x"52713370",x"81ff0652",x"5470802e",x"9d387233",x"5570752e",x"09810695",x"38811281",x"14713370",x"81ff0654",x"56545270",x"e5387233",x"557381ff",x"067581ff",x"06717131",x"880c5252",x"873d0d04",x"710970f7",x"fbfdff14",x"0670f884",x"82818006",x"51515170",x"97388414",x"84167108",x"54565471",x"75082edc",x"38737554",x"52ff9639",x"800b880c",x"873d0d04",x"ff3d0d9f",x"980bfc05",x"70085252",x"70ff2e91",x"38702dfc",x"12700852",x"5270ff2e",x"098106f1",x"38833d0d",x"0404eb83",x"3f040000",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"0000093d",x"0000096f",x"00000917",x"000007a2",x"000009c6",x"000009dd",x"00000835",x"000008c4",x"0000074e",x"000009f1",x"01090600",x"00006f80",x"05b8d800",x"b4010f00",x"00000000",x"00000000",x"00000000",x"00000fa0",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
